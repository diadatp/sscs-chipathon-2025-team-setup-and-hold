* NGSPICE file created from gf180mcu_sah_sc_aoi222_1.ext - technology: gf180mcuD

.subckt gf180mcu_sah_sc_aoi222_1 VSS VDD Y A1 A2 B1 B2 C2 C1
X0 VDD.t1 A2.t0 a_n3268_1558# VDD.t0 pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1 a_n3268_1558# B1.t0 a_n2938_1558# VDD.t3 pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X2 VSS.t2 C2.t0 a_n2412_658# VSS.t1 nfet_03v3 ad=0.425p pd=2.7u as=0.102p ps=1.09u w=0.85u l=0.3u
X3 a_n2412_658# C1.t0 Y.t3 VSS.t8 nfet_03v3 ad=0.102p pd=1.09u as=0.425p ps=2.7u w=0.85u l=0.3u
X4 Y.t4 C1.t1 a_n2938_1558# VDD.t7 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 a_n3268_1558# A1.t0 VDD.t6 VDD.t5 pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X6 Y.t0 A2.t1 a_n3268_658# VSS.t0 nfet_03v3 ad=0.425p pd=2.7u as=0.102p ps=1.09u w=0.85u l=0.3u
X7 a_n2938_1558# C2.t1 Y.t1 VDD.t2 pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X8 a_n3268_658# A1.t1 VSS.t4 VSS.t3 nfet_03v3 ad=0.102p pd=1.09u as=0.425p ps=2.7u w=0.85u l=0.3u
X9 a_n2938_1558# B2.t0 a_n3268_1558# VDD.t4 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X10 Y.t2 B2.t1 a_n2840_658# VSS.t5 nfet_03v3 ad=0.425p pd=2.7u as=0.102p ps=1.09u w=0.85u l=0.3u
X11 a_n2840_658# B1.t1 VSS.t7 VSS.t6 nfet_03v3 ad=0.102p pd=1.09u as=0.425p ps=2.7u w=0.85u l=0.3u
R0 A2.n0 A2.t1 63.1455
R1 A2.n0 A2.t0 54.5072
R2 A2 A2.n0 12.5106
R3 VDD.n7 VDD.t0 345.312
R4 VDD.t4 VDD.t7 265.625
R5 VDD.n6 VDD.t5 239.062
R6 VDD.t3 VDD.n3 217.189
R7 VDD.n2 VDD.t2 207.812
R8 VDD.n7 VDD.t3 154.689
R9 VDD.n4 VDD.t5 145.413
R10 VDD.t7 VDD.n2 57.813
R11 VDD.n3 VDD.t4 48.438
R12 VDD.t0 VDD.n6 26.563
R13 VDD.n2 VDD.n0 12.7535
R14 VDD.n3 VDD.n0 12.6005
R15 VDD.n8 VDD.n7 12.6005
R16 VDD.n6 VDD.n5 12.6005
R17 VDD.n4 VDD.t6 3.29819
R18 VDD.n1 VDD.t1 3.29819
R19 VDD.n5 VDD.n4 0.1535
R20 VDD.n8 VDD.n1 0.0879286
R21 VDD VDD.n0 0.0834286
R22 VDD VDD.n8 0.0705714
R23 VDD.n5 VDD.n1 0.0660714
R24 B1.n0 B1.t0 71.0538
R25 B1.n0 B1.t1 42.7075
R26 B1 B1.n0 12.5151
R27 C2.n0 C2.t1 70.2044
R28 C2.n0 C2.t0 42.5252
R29 C2 C2.n0 12.514
R30 VSS.n8 VSS.n7 758.333
R31 VSS.n4 VSS.t8 723.284
R32 VSS.t6 VSS.t5 344.118
R33 VSS.t3 VSS.t0 344.118
R34 VSS.n3 VSS.t1 309.07
R35 VSS.t5 VSS.n4 296.324
R36 VSS.n5 VSS.t3 281.233
R37 VSS.n7 VSS.t0 143.382
R38 VSS.n8 VSS.t6 117.892
R39 VSS.t8 VSS.n3 35.0495
R40 VSS.n3 VSS.n2 10.4005
R41 VSS.n4 VSS.n0 10.4005
R42 VSS.n9 VSS.n8 10.4005
R43 VSS.n7 VSS.n6 10.4005
R44 VSS.n2 VSS.t2 8.73474
R45 VSS.n5 VSS.t4 8.61774
R46 VSS.n1 VSS.t7 8.61774
R47 VSS.n2 VSS.n0 0.1535
R48 VSS.n6 VSS.n5 0.1535
R49 VSS.n6 VSS.n1 0.122643
R50 VSS VSS.n0 0.0834286
R51 VSS VSS.n9 0.0705714
R52 VSS.n9 VSS.n1 0.0313571
R53 C1.n0 C1.t0 59.6523
R54 C1.n0 C1.t1 53.4643
R55 C1 C1.n0 12.5106
R56 Y.n1 Y.t0 9.3555
R57 Y.n1 Y.t2 8.61594
R58 Y.n2 Y.t3 8.61594
R59 Y Y.n0 6.69811
R60 Y Y.n2 5.62461
R61 Y.n0 Y.t1 1.13285
R62 Y.n0 Y.t4 1.13285
R63 Y.n2 Y.n1 0.196152
R64 A1.n0 A1.t1 78.8725
R65 A1.n0 A1.t0 37.3842
R66 A1 A1.n0 12.5162
R67 B2.n0 B2.t0 86.6272
R68 B2.n0 B2.t1 36.0618
R69 B2 B2.n0 12.5151
C0 a_n3268_1558# Y 0.00435f
C1 B1 a_n2938_1558# 0.0566f
C2 C2 C1 0.12067f
C3 A1 C1 0
C4 C2 A2 0
C5 B2 C1 0.1032f
C6 A1 A2 0.1265f
C7 B1 VDD 0.09421f
C8 a_n3268_658# Y 0.00307f
C9 B2 A2 0.00238f
C10 B1 a_n3268_1558# 0.03133f
C11 C1 Y 0.15824f
C12 VDD a_n2938_1558# 0.39059f
C13 a_n2938_1558# a_n3268_1558# 0.36504f
C14 A2 Y 0.03334f
C15 VDD a_n3268_1558# 0.41968f
C16 B1 C1 0.00408f
C17 C1 a_n2938_1558# 0.07022f
C18 B1 A2 0.04403f
C19 Y a_n2840_658# 0.006f
C20 A2 a_n2938_1558# 0.00275f
C21 C2 A1 0
C22 C2 B2 0.00154f
C23 VDD a_n3268_658# 0
C24 A1 B2 0.00149f
C25 a_n3268_658# a_n3268_1558# 0
C26 C1 VDD 0.08828f
C27 C1 a_n3268_1558# 0
C28 C2 Y 0.12416f
C29 VDD A2 0.11846f
C30 B1 a_n2840_658# 0.00116f
C31 A1 Y 0.01468f
C32 A2 a_n3268_1558# 0.03397f
C33 B2 Y 0.16178f
C34 C2 B1 0.00744f
C35 A1 B1 0.00229f
C36 C2 a_n2938_1558# 0.059f
C37 C1 A2 0.0125f
C38 B1 B2 0.12682f
C39 A1 a_n2938_1558# 0
C40 B2 a_n2938_1558# 0.05309f
C41 B1 Y 0.06556f
C42 a_n2938_1558# Y 0.45803f
C43 C2 VDD 0.09158f
C44 A1 VDD 0.12957f
C45 C2 a_n3268_1558# 0
C46 A1 a_n3268_1558# 0.01493f
C47 B2 VDD 0.08581f
C48 Y a_n2412_658# 0.00675f
C49 B2 a_n3268_1558# 0.01611f
C50 VDD Y 0.06673f
C51 Y VSS 0.79808f
C52 C2 VSS 0.62196f
C53 C1 VSS 0.49701f
C54 B2 VSS 0.5476f
C55 B1 VSS 0.53489f
C56 A2 VSS 0.54208f
C57 A1 VSS 0.57838f
C58 VDD VSS 3.09588f
C59 a_n2412_658# VSS 0.00586f
C60 a_n2840_658# VSS 0.00586f
C61 a_n3268_658# VSS 0.00586f
C62 a_n2938_1558# VSS 0.12889f
C63 a_n3268_1558# VSS 0.12917f
.ends

